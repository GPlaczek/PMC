library IEEE;
	use IEEE.std_logic_1164.all;
	
entity counter is
	port (bus_in: in std_logic_vector(7 downto 0));
end entity;

architecture empty of counter is
begin
end architecture;
